library ieee;
use ieee.std_logic_1164.all;
use ieee.math_real.all; 



package my_package is
	type my_arr_bit is array (0 to 4) of std_logic_vector(7 downto 0);	 
	type my_arr_int is array (0 to 4) of integer;
end my_package;	 

	