library ieee;
use ieee.std_logic_1164.all;
use ieee.math_real.all; 



package my_arr is
	type arr is array (0 to 7) of integer;
end my_arr;	 