library ieee;
use ieee.std_logic_1164.all;
use ieee.math_real.all; 



package my_package is
	type matrix is array (0 to 2, 0 to 2) of std_logic_vector(3 downto 0);
end my_package;	 

	